module dff(
  output reg Q,
  input D,
  input Clk)
  
endmodule
